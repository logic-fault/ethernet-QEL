** Profile: "SCHEMATIC1-SIM_MAIN"  [ H:\ETHERNET-QEL\SIMULATION\QEL_Drive\qel_drive-SCHEMATIC1-SIM_MAIN.sim ] 

** Creating circuit file "qel_drive-SCHEMATIC1-SIM_MAIN.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10s 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\qel_drive-SCHEMATIC1.net" 


.END
